library ieee;
use ieee.std_logic_1164.all;

entity FlipFlopD is
	port( 
			clock: in std_logic;
			reset: in std_logic;
			D: in std_logic;
	      Q: out std_logic
	    );
end FlipFlopD;

architecture RTL of FlipFlopD is
begin
	process(clock, reset)
	begin
		if (reset = '1') then
			Q <= '0';
		elsif (clock = '1' and clock'event) then
			Q <= D;
		end if;
	end process;
end RTL;